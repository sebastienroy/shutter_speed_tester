.title KiCad schematic
H3 MountingHole
H2 MountingHole
H1 MountingHole
H4 MountingHole
J4 Net-_A1-Pad30_ GND Power
A1 NC_01 NC_02 NC_03 GND Net-_A1-Pad5_ Net-_A1-Pad6_ Net-_A1-Pad7_ Net-_A1-Pad8_ NC_04 NC_05 NC_06 NC_07 NC_08 NC_09 NC_10 NC_11 NC_12 NC_13 NC_14 NC_15 NC_16 NC_17 Net-_A1-Pad23_ Net-_A1-Pad24_ NC_18 NC_19 Net-_A1-Pad27_ NC_20 GND Net-_A1-Pad30_ Arduino_Nano_v3.x
R1 Net-_A1-Pad5_ GND 1meg
J3 GND Net-_A1-Pad27_ Net-_A1-Pad23_ Net-_A1-Pad24_ LCD
Q1 GND Net-_Q1-Pad2_ Net-_Q1-Pad3_ PN2222A
R4 Net-_A1-Pad6_ Net-_Q1-Pad2_ 1k
R2 Net-_J2-Pad1_ Net-_Q1-Pad3_ 220
SW1 Net-_A1-Pad7_ Net-_A1-Pad27_ Reset switch
R3 Net-_A1-Pad7_ GND 10k
D1 Net-_D1-Pad1_ Net-_A1-Pad8_ Control LED
R5 Net-_D1-Pad1_ GND 1k
J2 Net-_J2-Pad1_ Net-_A1-Pad27_ Light source LED
J1 Net-_A1-Pad5_ Net-_A1-Pad27_ Light Sensor
.end
